----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:41:26 05/08/2012 
-- Design Name: 
-- Module Name:    ADC_data_handler_v3 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;

use work.ADC_data_handler_package.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ADC_data_handler_v4 is

  port (
    reset : in std_logic;
    clk   : in std_logic;

    testmode_rst : in std_logic;
    testmode_col : in std_logic;

    start_of_img : in std_logic;  -- this signal is generated by the user (using the sequencer) and has to arrive before the first trigger
    end_of_img   : in std_logic;  -- this signal is generated by the user (using the sequencer) and has to arrive after the last  ADC trasfer
    end_sequence : in std_logic;  -- this signal is the end of sequence generated by the sequencer and is used as a timeot to generate EOF.

    trigger : in std_logic;  -- this signal start the operations (ADC conv and send data to PGP)
--              image_size                      : in  std_logic_vector(31 downto 0);    -- this is the image size 
--              en_load_image_size      : in  std_logic;                                                                -- load the image size into register

    en_test_mode : in std_logic;  -- register enable for pattern test mode
    test_mode_in : in std_logic;        -- test mode in 

    en_load_ccd_sel : in  std_logic;    -- register enable for CCD enable
    ccd_sel_in      : in  std_logic_vector(2 downto 0);  -- register to select which CCD acquire (1, 2 or 3) 
    ccd_sel_out     : out std_logic_vector(2 downto 0);  -- register to select which CCD acquire (1, 2 or 3) 

    SOT          : out std_logic;       -- Start of Image
    EOT          : out std_logic;       -- End of Image
    write_enable : out std_logic;       -- signal to write the image in the PGP

    test_mode_enb_out : out std_logic;
--              image_size_out                  : out std_logic_vector(31 downto 0);    -- Image size read (for RCE)


    data_out : out std_logic_vector(17 downto 0);  -- 18 bits ADC word 

    adc_data_ccd_1 : in  std_logic_vector(15 downto 0);  -- CCD ADC data 
    adc_cnv_ccd_1  : out std_logic;                      -- ADC conv
    adc_sck_ccd_1  : out std_logic;                      -- ADC serial clock

    adc_data_ccd_2 : in  std_logic_vector(15 downto 0);  -- CCD ADC data 
    adc_cnv_ccd_2  : out std_logic;                      -- ADC conv
    adc_sck_ccd_2  : out std_logic;                      -- ADC serial clock

    adc_data_ccd_3 : in  std_logic_vector(15 downto 0);  -- CCD ADC data 
    adc_cnv_ccd_3  : out std_logic;                      -- ADC conv
    adc_sck_ccd_3  : out std_logic                       -- ADC serial clock

    );

end ADC_data_handler_v4;

architecture Behavioral of ADC_data_handler_v4 is


  component ADC_data_handler_fsm_v4 is
    port (
      reset        : in  std_logic;
      clk          : in  std_logic;
      trigger      : in  std_logic;
--       cnt_end                  : in  std_logic;
      start_of_img : in  std_logic;  -- this signal is generated by the user (using the sequencer) and has to arrive before the first trigger
      end_of_img   : in  std_logic;  -- this signal is generated by the user (using the sequencer) and has to arrive after the last  ADC trasfer
      end_sequence : in  std_logic;  -- this signal is the end of sequence generated by the sequencer and is used as a timeot to generate EOF.
      ccd_sel      : in  std_logic_vector(2 downto 0);
      data_ccd_1   : in  array1618;
      data_ccd_2   : in  array1618;
      data_ccd_3   : in  array1618;
      cnt_en       : out std_logic;
      init_cnt     : out std_logic;
      SOT          : out std_logic;
      EOT          : out std_logic;
      write_enable : out std_logic;
      handler_busy : out std_logic;
      data_out     : out std_logic_vector(17 downto 0)
      );
  end component;

  component generic_counter_comparator_ce_init is
    generic (length_cnt : integer);
    port (
      reset     : in  std_logic;        -- syncronus reset
      clk       : in  std_logic;        -- clock
      max_value : in  std_logic_vector (length_cnt downto 0);  -- maximum value the counter has to count
      enable    : in  std_logic;        -- enable
      init      : in  std_logic;
      cnt_end   : out std_logic;  -- signal = 1 when the counter reach the maximum
      q_out     : out std_logic_vector(length_cnt downto 0));
  end component;

  component generic_reg_ce_init is
    generic (width : integer);
    port (
      reset    : in  std_logic;         -- syncronus reset
      clk      : in  std_logic;         -- clock
      ce       : in  std_logic;         -- clock enable
      init     : in  std_logic;  -- signal to reset the reg (active high)
      data_in  : in  std_logic_vector(width downto 0);   -- data in
      data_out : out std_logic_vector(width downto 0));  -- data out
  end component;

  component generic_reg_ce_init_1 is
    generic (width : integer);
    port (
      reset    : in  std_logic;         -- syncronus reset
      clk      : in  std_logic;         -- clock
      ce       : in  std_logic;         -- clock enable
      init     : in  std_logic;  -- signal to reset the reg (active high)
      data_in  : in  std_logic_vector(width downto 0);   -- data in
      data_out : out std_logic_vector(width downto 0));  -- data out
  end component;

  component readadcs_v5 is
    generic (
      conv_time        : integer := 50;
      sclk_half_period : integer := 1;
      test_time        : integer := 500;
      col_incr_val     : integer := 10;
      pix_incr_val     : integer := 8
      );
    port(
      clk          : in  std_logic;
      reset        : in  std_logic;
      start_conv   : in  std_logic;
      testmode_enb : in  std_logic;
      testmode_rst : in  std_logic;
      testmode_col : in  std_logic;
      adc_data     : in  std_logic_vector(15 downto 0);
      adc_cnv      : out std_logic;
      adc_sck      : out std_logic;
      data_ready   : out std_logic;
      adc_ch       : out array1618

      );
  end component;

  component ff_ce is
    port (

      reset : in std_logic;

      clk     : in std_logic;
      data_in : in std_logic;
      ce      : in std_logic;

      data_out : out std_logic); 
  end component;



  signal cnt_en   : std_logic;
--signal cnt_end                                : std_logic;
  signal init_cnt : std_logic;
--signal image_size_out_int             : std_logic_vector(31 downto 0);

  signal testmode_enb : std_logic;

  signal data_ready       : std_logic;
  signal data_ready_ccd_1 : std_logic;
  signal data_ready_ccd_2 : std_logic;
  signal data_ready_ccd_3 : std_logic;

  signal trigger_ccd_1 : std_logic;
  signal trigger_ccd_2 : std_logic;
  signal trigger_ccd_3 : std_logic;

  signal end_sequence_stretch     : std_logic;
  signal end_sequence_stretch_inv : std_logic;
  signal handler_busy             : std_logic;
  signal stretch_reset            : std_logic;

  signal ADC_CCD_1 : array1618;
  signal ADC_CCD_2 : array1618;
  signal ADC_CCD_3 : array1618;

  signal ccd_sel : std_logic_vector(2 downto 0);

begin


  test_mode_enb_out <= testmode_enb;
--      image_size_out          <= image_size_out_int;

  trigger_ccd_1 <= trigger and ccd_sel(0);
  trigger_ccd_2 <= trigger and ccd_sel(1);
  trigger_ccd_3 <= trigger and ccd_sel(2);

  data_ready <= data_ready_ccd_1 or data_ready_ccd_2 or data_ready_ccd_3;

  ccd_sel_out <= ccd_sel;

  stretch_reset            <= reset or (not handler_busy);
  end_sequence_stretch_inv <= not end_sequence_stretch;

  ADC_data_handler_fsm_v4_0 : ADC_data_handler_fsm_v4
    port map (
      reset        => reset,
      clk          => clk,
      trigger      => data_ready,
--      cnt_end          => cnt_end,
      start_of_img => start_of_img,
      end_of_img   => end_of_img,
      end_sequence => end_sequence_stretch,
      ccd_sel      => ccd_sel,
      data_ccd_1   => ADC_CCD_1,
      data_ccd_2   => ADC_CCD_2,
      data_ccd_3   => ADC_CCD_3,
      cnt_en       => cnt_en,
      init_cnt     => init_cnt,
      SOT          => SOT,
      EOT          => EOT,
      write_enable => write_enable,
      handler_busy => handler_busy,
      data_out     => data_out
      );


  end_seq_stretch : ff_ce
    port map (
      reset    => stretch_reset,
      clk      => clk,
      data_in  => end_sequence,
      ce       => end_sequence_stretch_inv,
      data_out => end_sequence_stretch
      ); 

  sel_ccd_reg : generic_reg_ce_init_1
    generic map (
      width => 2)
    port map(
      reset    => reset,
      clk      => clk,
      ce       => en_load_ccd_sel,
      init     => '0',
      data_in  => ccd_sel_in,
      data_out => ccd_sel);


  trigger_counter : generic_counter_comparator_ce_init
    generic map (
      length_cnt => 31)
    port map(
      reset     => reset,
      clk       => clk,
      max_value => x"00000000",
      enable    => cnt_en,
      init      => init_cnt,
      cnt_end   => open,
      q_out     => open);
--
--
--  trigger_counter_reg : generic_reg_ce_init
--    generic map (
--      width    => 31)
--    port map(
--      reset    => reset,
--      clk      => clk,
--      ce       => en_load_image_size,
--      init     => '0',
--      data_in  => image_size,
--      data_out => image_size_out_int);

  readadcs_v5_0_ccd1 : readadcs_v5
    generic map (
      conv_time        => 75,
      sclk_half_period => 2,
      test_time        => 150,
      col_incr_val     => 10,
      pix_incr_val     => 8
      )
    port map(
      clk          => clk,
      reset        => reset,
      start_conv   => trigger_ccd_1,
      testmode_enb => testmode_enb,
      testmode_rst => testmode_rst,
      testmode_col => testmode_col,
      adc_data     => adc_data_ccd_1,
      adc_cnv      => adc_cnv_ccd_1,
      adc_sck      => adc_sck_ccd_1,
      data_ready   => data_ready_ccd_1,
      adc_ch       => ADC_CCD_1
      );

  readadcs_v5_0_ccd2 : readadcs_v5
    generic map (
      conv_time        => 75,
      sclk_half_period => 2,
      test_time        => 150,
      col_incr_val     => 10,
      pix_incr_val     => 8
      )
    port map(
      clk          => clk,
      reset        => reset,
      start_conv   => trigger_ccd_2,
      testmode_enb => testmode_enb,
      testmode_rst => testmode_rst,
      testmode_col => testmode_col,
      adc_data     => adc_data_ccd_2,
      adc_cnv      => adc_cnv_ccd_2,
      adc_sck      => adc_sck_ccd_2,
      data_ready   => data_ready_ccd_2,
      adc_ch       => ADC_CCD_2
      );

  readadcs_v5_0_ccd3 : readadcs_v5
    generic map (
      conv_time        => 75,
      sclk_half_period => 2,
      test_time        => 150,
      col_incr_val     => 10,
      pix_incr_val     => 8
      )
    port map(
      clk          => clk,
      reset        => reset,
      start_conv   => trigger_ccd_3,
      testmode_enb => testmode_enb,
      testmode_rst => testmode_rst,
      testmode_col => testmode_col,
      adc_data     => adc_data_ccd_3,
      adc_cnv      => adc_cnv_ccd_3,
      adc_sck      => adc_sck_ccd_3,
      data_ready   => data_ready_ccd_3,
      adc_ch       => ADC_CCD_3
      );

  test_mode_ff : ff_ce
    port map (

      reset => reset,

      clk     => clk,
      data_in => test_mode_in,
      ce      => en_test_mode,

      data_out => testmode_enb
      ); 

end Behavioral;

